module DataMemory #(
    parameter integer MEM_DEPTH = 16384
) (
    input         reset,
    input         clk,
    input  [31:0] addr,       // address of the data memory
    input  [31:0] din,        // data to be written
    input         mem_read,   // is read signal driven?
    input         mem_write,  // is write signal driven?
    output [31:0] dout        // output of the data memory at addr
);
  integer i;
  // Data memory
  reg [31:0] mem[MEM_DEPTH];
  // Do not touch dmem_addr
  wire [31:0] dmem_addr;
  assign dmem_addr = {addr >> 2};

  // Asynchrnously read data from the memory
  // Synchronously write data to the memory
  assign dout = (mem_read) ? mem[dmem_addr] : 32'b0;
  always @(posedge clk) begin
    if (reset) begin
      for (i = 0; i < MEM_DEPTH; i = i + 1)
      // DO NOT TOUCH COMMENT BELOW
      /* verilator lint_off BLKSEQ */
      mem[i] = 32'b0;
      /* verilator lint_on BLKSEQ */
      // DO NOT TOUCH COMMENT ABOVE
    end else begin
      if (mem_write) mem[dmem_addr] <= din;
    end
  end
endmodule


